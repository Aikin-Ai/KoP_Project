library ieee;
use ieee.std_logic_1164.all;

entity button_controller is

	port 
	(
		clk		  : in std_logic;
		button_in  : in std_logic;
		button_out : out std_logic
	);

end button_controller;

architecture rtl of button_controller is

begin

	

end rtl;
